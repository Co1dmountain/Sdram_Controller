module Sdram_write(
		// input
);












endmodule