module uart_tx(
		//system signals
		input					sclk				,
		input					s_rst_n				,
		//tx_flag
		input					tx_flag				,
		//UART Interface
		output					rs232_tx			,
		//others
		output	reg		[7:0]	tx_data				,

);

	//define parameter and internal signals
	
	//main code
	
	

	

	
	
	
	
	
	
	
	
	
	
	
endmodule