module Sdram_write(
		// input
		input 				sys_clk					,
		input				sys_rst_n				,
		// write_en?
		input				write_en				,
		
		// output
		output				write_req				,
		output				write_end
);

	//// define ////
	// 定义指令、计数器、寄存器、状态机状态（写数据过程的状态机，
	// 在顶层文件中应该还有写状态这一状态，当顶层状态机进入写数据状态，
	// 就进入该模块进行写数据操作）
	
	
	
	//// main code ////
	
	
	
	
	
	
	
	
	


endmodule